`timescale 1ns / 1ps

module test_sum;
    reg clk = 0;
    reg rst = 0;
    
    // ������ ����������
    wire [15:0] ACC;
    wire halted;
    
    // ��������� ��������� �������
    always #1 clk <= ~clk;
    
    // ��������� ����������
    cpu dut(
        .clk(clk),
        .rst(rst),
        .ACC(ACC),
        .halted(halted)
    );
    
endmodule